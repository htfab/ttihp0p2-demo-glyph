`ifndef DIV3_ROM_H
`define DIV3_ROM_H

// Division-by-3 lookup table

module div3_rom(
    input wire [6:0] in,
    output wire [5:0] out
);
	reg [5:0] d[0:119];
	assign out = d[in];
	initial begin
		d[  0] = 6'd0;
		d[  1] = 6'd0;
		d[  2] = 6'd0;
		d[  3] = 6'd1;
		d[  4] = 6'd1;
		d[  5] = 6'd1;
		d[  6] = 6'd2;
		d[  7] = 6'd2;
		d[  8] = 6'd2;
		d[  9] = 6'd3;
		d[ 10] = 6'd3;
		d[ 11] = 6'd3;
		d[ 12] = 6'd4;
		d[ 13] = 6'd4;
		d[ 14] = 6'd4;
		d[ 15] = 6'd5;
		d[ 16] = 6'd5;
		d[ 17] = 6'd5;
		d[ 18] = 6'd6;
		d[ 19] = 6'd6;
		d[ 20] = 6'd6;
		d[ 21] = 6'd7;
		d[ 22] = 6'd7;
		d[ 23] = 6'd7;
		d[ 24] = 6'd8;
		d[ 25] = 6'd8;
		d[ 26] = 6'd8;
		d[ 27] = 6'd9;
		d[ 28] = 6'd9;
		d[ 29] = 6'd9;
		d[ 30] = 6'd10;
		d[ 31] = 6'd10;
		d[ 32] = 6'd10;
		d[ 33] = 6'd11;
		d[ 34] = 6'd11;
		d[ 35] = 6'd11;
		d[ 36] = 6'd12;
		d[ 37] = 6'd12;
		d[ 38] = 6'd12;
		d[ 39] = 6'd13;
		d[ 40] = 6'd13;
		d[ 41] = 6'd13;
		d[ 42] = 6'd14;
		d[ 43] = 6'd14;
		d[ 44] = 6'd14;
		d[ 45] = 6'd15;
		d[ 46] = 6'd15;
		d[ 47] = 6'd15;
		d[ 48] = 6'd16;
		d[ 49] = 6'd16;
		d[ 50] = 6'd16;
		d[ 51] = 6'd17;
		d[ 52] = 6'd17;
		d[ 53] = 6'd17;
		d[ 54] = 6'd18;
		d[ 55] = 6'd18;
		d[ 56] = 6'd18;
		d[ 57] = 6'd19;
		d[ 58] = 6'd19;
		d[ 59] = 6'd19;
		d[ 60] = 6'd20;
		d[ 61] = 6'd20;
		d[ 62] = 6'd20;
		d[ 63] = 6'd21;
		d[ 64] = 6'd21;
		d[ 65] = 6'd21;
		d[ 66] = 6'd22;
		d[ 67] = 6'd22;
		d[ 68] = 6'd22;
		d[ 69] = 6'd23;
		d[ 70] = 6'd23;
		d[ 71] = 6'd23;
		d[ 72] = 6'd24;
		d[ 73] = 6'd24;
		d[ 74] = 6'd24;
		d[ 75] = 6'd25;
		d[ 76] = 6'd25;
		d[ 77] = 6'd25;
		d[ 78] = 6'd26;
		d[ 79] = 6'd26;
		d[ 80] = 6'd26;
		d[ 81] = 6'd27;
		d[ 82] = 6'd27;
		d[ 83] = 6'd27;
		d[ 84] = 6'd28;
		d[ 85] = 6'd28;
		d[ 86] = 6'd28;
		d[ 87] = 6'd29;
		d[ 88] = 6'd29;
		d[ 89] = 6'd29;
		d[ 90] = 6'd30;
		d[ 91] = 6'd30;
		d[ 92] = 6'd30;
		d[ 93] = 6'd31;
		d[ 94] = 6'd31;
		d[ 95] = 6'd31;
		d[ 96] = 6'd32;
		d[ 97] = 6'd32;
		d[ 98] = 6'd32;
		d[ 99] = 6'd33;
		d[100] = 6'd33;
		d[101] = 6'd33;
		d[102] = 6'd34;
		d[103] = 6'd34;
		d[104] = 6'd34;
		d[105] = 6'd35;
		d[106] = 6'd35;
		d[107] = 6'd35;
		d[108] = 6'd36;
		d[109] = 6'd36;
		d[110] = 6'd36;
		d[111] = 6'd37;
		d[112] = 6'd37;
		d[113] = 6'd37;
		d[114] = 6'd38;
		d[115] = 6'd38;
		d[116] = 6'd38;
		d[117] = 6'd39;
		d[118] = 6'd39;
		d[119] = 6'd39;
	end

endmodule

`endif
